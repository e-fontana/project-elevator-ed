module block_doors;
endmodule