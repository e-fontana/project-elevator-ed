module frequency_door #(parameter door_time = 2) (clk, move_handler, door_clk);
	input clk, move_handler;
	output reg door_clk;

	reg [25:0] counter = 0;

	always @(posedge move_handler) begin
		counter <= 0;
	end
	
	always @(posedge clk) begin
		if (counter < door_time) begin
			counter <= counter + 1;
			door_clk <= 1'b0;
		end else begin
			counter <= 1'b0;
			door_clk <= ~door_clk;
		end
	end
endmodule