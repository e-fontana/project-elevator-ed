module moviment_direction_tb;
    
endmodule