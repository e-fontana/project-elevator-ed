`include "./emergency/design.v"

module emergency_tb;
    
endmodule