module moviment_direction;
    
endmodule