module door_block_tb;
    
endmodule