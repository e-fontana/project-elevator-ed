module door_status;
endmodule