module tb;
endmodule