`include "frequency_divisor.v"

`include "click_handler/location.v"

`include "emergency/sos_handler.v"
`include "emergency/door_situation.v"
`include "emergency/weight_control.v"

`include "position/queue.v"
`include "position/moviment.v"

module TOP(clk);
    input clk;

endmodule