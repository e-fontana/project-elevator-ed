module door_block;
    
endmodule