module moviment_authorization;
    
endmodule