module moviment_authorization_tb;
    
endmodule