module led_disable(goal_floor, led1, led2, led3);
endmodule