module weight_control_tb;
endmodule